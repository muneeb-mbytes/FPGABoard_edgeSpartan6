dgdddg
